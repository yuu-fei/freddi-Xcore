///////////////////////////////////////////////////////////////////////////////
//
// Copyright Freddi, UESTC 
//
///////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps
//-----------------------------------------------------------------------------
//
// Project    : Xcore fifo
// File       : Xcore_fifo.v
// Module     : Xcore_fifo.v(sync fifo)
// Author     : Yufei Fu(fuyufei083X@gmail.com)
// Date       : 2022-9-29
// Version    : v1.0
// Description: sync fifo with data valid flag
//
// ----------------------------------------------------------------------------


module Xcore_fifo #(
	parameter DW = 8
)(
	input sys_clk,
	input sys_rst,

);


endmodule
