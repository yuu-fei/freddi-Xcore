///////////////////////////////////////////////////////////////////////////////
//
// Copyright Freddi, UESTC 
//
///////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps
//-----------------------------------------------------------------------------
//
// Project    : Xcore regfile module in id section
// File       : Xcore_id_regf.v
// Module     : Xcore_id_regf.v(regfile)
// Author     : Yufei Fu(fuyufei083X@gmail.com)
// Date       : 2022-9-25
// Version    : v1.0
// Description: Regfile to hold using data 
//				bypass input is considered
//				two points;
//              register x0 is always 0
//              read is asynchronous while write shoulld be synchronous
//              use macro to selectively activate BYPASS datapath
//              
// ----------------------------------------------------------------------------
`include "./rtl/include/params.v"
module Xcore_id_regf(
	input			regf_clk,
	input			regf_rst,
	input			regwrite, // 0 is read while 1 is write
	//adress input
	input [4:0]		instr_id_rs1,
	input [4:0]		instr_id_rs2,
	input [4:0]		id_wd,

	//data input & output
	input [`WIDTH]	id_write_data,
	output [`WIDTH] id_read_data1,
	output [`WIDTH] id_read_data2

);
wire [`WIDTH]	 en; //this enable signal may be generated by outward control module
wire [`WIDTH]	 gpr_r[31:0];
//set regfile 32*32 using general dfflr

genvar i;

generate 
	for(i=0;i<32;i=i+1) begin: generate_regfile
		if(i==0) begin: is_x0
			assign en[i] = 'd0;
			assign gpr_r[i] = 'd0;
			Xcore_gnrl_dfflr #(32) dfflr_gp(regf_clk, en[i], regf_rst, id_write_data, gpr_r[i]);
		end
		else begin
			assign en[i] = regwrite&(id_wd==i);
			Xcore_gnrl_dfflr #(32) dfflr_gp(regf_clk, en[i], regf_rst, id_write_data, gpr_r[i]);
		end
	end
endgenerate

`ifdef XCORE_HAS_BYPASS
	// wriet-data when conflict at the same time
	assign 	id_read_data1 = (regwrite&(id_wd==instr_id_rs1)&(instr_id_rs1!=0)) ? id_write_data : gpr_r[instr_id_rs1];
	assign	id_read_data2 = (regwrite&(id_wd==instr_id_rs2)&(instr_id_rs2!=0)) ? id_write_data : gpr_r[instr_id_rs2];
`else
	assign id_read_data1 = gpr_r[instr_id_rs1];
	assign id_read_data2 = gpr_r[instr_id_rs2];
`endif
endmodule

